`timescale 1ps / 1ps
`default_nettype none
